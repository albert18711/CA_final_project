module ALUControl (
	IR_func,
	ALUOp,
	Jr_sel,
	ALUctrl
);

	input [5:0] IR_func;
	input [1:0] ALUOp;
	output reg Jr_sel;
	output reg [3:0] ALUctrl;



endmodule